LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

package generated is

  function builtin_rom(addr : in std_logic_vector(15 downto 1)) return std_logic_vector;

end package;

package body generated is

  function builtin_rom(addr : in std_logic_vector(15 downto 1)) return std_logic_vector is
  begin
    case to_integer(unsigned(addr & "0")) is
      when 16#0000# => return "0000001000001000";
      when 16#0002# => return "0000000000001010";
      when 16#0004# => return "0000000110100000";
      when 16#0006# => return "0000000101111110";
      when 16#0008# => return "0000000111000110";
      when 16#000A# => return "0011110000001000";
      when 16#000C# => return "0110000100000000";
      when 16#000E# => return "0000000100001000";
      when 16#0010# => return "0000000000100000";
      when 16#0012# => return "0000010100001000";
      when 16#0014# => return "0000000000000010";
      when 16#0016# => return "0000001000001000";
      when 16#0018# => return "0000000101111110";
      when 16#001A# => return "0000000000011000";
      when 16#001C# => return "0000001000001000";
      when 16#001E# => return "0000000010000100";
      when 16#0020# => return "0101101100011011";
      when 16#0022# => return "0001101101001000";
      when 16#0024# => return "0100101001011011";
      when 16#0026# => return "0011110100101110";
      when 16#0028# => return "0011110100111101";
      when 16#002A# => return "0011110100111101";
      when 16#002C# => return "0011110100111101";
      when 16#002E# => return "0011110100111101";
      when 16#0030# => return "0011110100111101";
      when 16#0032# => return "0011110100111101";
      when 16#0034# => return "0011110100111101";
      when 16#0036# => return "0011110100111101";
      when 16#0038# => return "0011110100111101";
      when 16#003A# => return "0011110100111101";
      when 16#003C# => return "0011110100111101";
      when 16#003E# => return "0011110100111101";
      when 16#0040# => return "0010111000111101";
      when 16#0042# => return "0000101000001101";
      when 16#0044# => return "0010000001111100";
      when 16#0046# => return "0101001101000001";
      when 16#0048# => return "0100010101001000";
      when 16#004A# => return "0010000001010100";
      when 16#004C# => return "0100111101001000";
      when 16#004E# => return "0100010101001101";
      when 16#0050# => return "0100001100100000";
      when 16#0052# => return "0100110101001111";
      when 16#0054# => return "0101010101010000";
      when 16#0056# => return "0100010101010100";
      when 16#0058# => return "0010000001010010";
      when 16#005A# => return "0100100101000010";
      when 16#005C# => return "0101001101001111";
      when 16#005E# => return "0111110000100000";
      when 16#0060# => return "0000101000001101";
      when 16#0062# => return "0011110100100111";
      when 16#0064# => return "0011110100111101";
      when 16#0066# => return "0011110100111101";
      when 16#0068# => return "0011110100111101";
      when 16#006A# => return "0011110100111101";
      when 16#006C# => return "0011110100111101";
      when 16#006E# => return "0011110100111101";
      when 16#0070# => return "0011110100111101";
      when 16#0072# => return "0011110100111101";
      when 16#0074# => return "0011110100111101";
      when 16#0076# => return "0011110100111101";
      when 16#0078# => return "0011110100111101";
      when 16#007A# => return "0011110100111101";
      when 16#007C# => return "0010011100111101";
      when 16#007E# => return "0000101000001101";
      when 16#0080# => return "0000101000001101";
      when 16#0084# => return "0001010000101000";
      when 16#0086# => return "0100000000000000";
      when 16#0088# => return "0000000000001101";
      when 16#008A# => return "0001010000101000";
      when 16#008C# => return "0100000000000000";
      when 16#008E# => return "0000000000111110";
      when 16#0090# => return "0001010000101000";
      when 16#0092# => return "0100000000000000";
      when 16#0094# => return "0000000000100000";
      when 16#0096# => return "0001010000101000";
      when 16#0098# => return "0100000000000000";
      when 16#009A# => return "0000000000100000";
      when 16#009C# => return "0001010000101000";
      when 16#009E# => return "0100000000000000";
      when 16#00A0# => return "0000000000001000";
      when 16#00A2# => return "0001110110001000";
      when 16#00A4# => return "0100000000000000";
      when 16#00A6# => return "0000001001101100";
      when 16#00A8# => return "0000000010100010";
      when 16#00AA# => return "0001010001001000";
      when 16#00AC# => return "0100000000000000";
      when 16#00AE# => return "0100010010110000";
      when 16#00B0# => return "0000000001101000";
      when 16#00B2# => return "0000001001101001";
      when 16#00B4# => return "0000000011000100";
      when 16#00B6# => return "0100010010110000";
      when 16#00B8# => return "0000000001100111";
      when 16#00BA# => return "0000001001101001";
      when 16#00BC# => return "0000000101101010";
      when 16#00BE# => return "0000000000011000";
      when 16#00C0# => return "0000001000001000";
      when 16#00C2# => return "0000000010000100";
      when 16#00C4# => return "0000000100001000";
      when 16#00C6# => return "0000000011010110";
      when 16#00C8# => return "0000010100001000";
      when 16#00CA# => return "0000000000000010";
      when 16#00CC# => return "0000001000001000";
      when 16#00CE# => return "0000000101111110";
      when 16#00D0# => return "0000000000011000";
      when 16#00D2# => return "0000001000001000";
      when 16#00D4# => return "0000000010000100";
      when 16#00D6# => return "0000101000001101";
      when 16#00D8# => return "0111011001100001";
      when 16#00DA# => return "0110100101100001";
      when 16#00DC# => return "0110000101101100";
      when 16#00DE# => return "0110110001100010";
      when 16#00E0# => return "0010000001100101";
      when 16#00E2# => return "0110111101100011";
      when 16#00E4# => return "0110110101101101";
      when 16#00E6# => return "0110111001100001";
      when 16#00E8# => return "0111001101100100";
      when 16#00EA# => return "0000110100111010";
      when 16#00EC# => return "0010000000001010";
      when 16#00EE# => return "0110100000100000";
      when 16#00F0# => return "0010000000100000";
      when 16#00F2# => return "0010000000101101";
      when 16#00F4# => return "0110100101100100";
      when 16#00F6# => return "0111000001110011";
      when 16#00F8# => return "0110000101101100";
      when 16#00FA# => return "0010000001111001";
      when 16#00FC# => return "0110010101101000";
      when 16#00FE# => return "0111000001101100";
      when 16#0100# => return "0000101000001101";
      when 16#0102# => return "0010000000100000";
      when 16#0104# => return "0110001001110010";
      when 16#0106# => return "0010110100100000";
      when 16#0108# => return "0111001000100000";
      when 16#010A# => return "0110000101100101";
      when 16#010C# => return "0010000001100100";
      when 16#010E# => return "0111100101100010";
      when 16#0110# => return "0110010101110100";
      when 16#0112# => return "0000101000001101";
      when 16#0114# => return "0010000000100000";
      when 16#0116# => return "0111011101110010";
      when 16#0118# => return "0010110100100000";
      when 16#011A# => return "0111001000100000";
      when 16#011C# => return "0110000101100101";
      when 16#011E# => return "0010000001100100";
      when 16#0120# => return "0110111101110111";
      when 16#0122# => return "0110010001110010";
      when 16#0124# => return "0000101000001101";
      when 16#0126# => return "0010000000100000";
      when 16#0128# => return "0110001001110111";
      when 16#012A# => return "0010110100100000";
      when 16#012C# => return "0111011100100000";
      when 16#012E# => return "0110100101110010";
      when 16#0130# => return "0110010101110100";
      when 16#0132# => return "0110001000100000";
      when 16#0134# => return "0111010001111001";
      when 16#0136# => return "0000110101100101";
      when 16#0138# => return "0010000000001010";
      when 16#013A# => return "0111011100100000";
      when 16#013C# => return "0010000001110111";
      when 16#013E# => return "0010000000101101";
      when 16#0140# => return "0111001001110111";
      when 16#0142# => return "0111010001101001";
      when 16#0144# => return "0010000001100101";
      when 16#0146# => return "0110111101110111";
      when 16#0148# => return "0110010001110010";
      when 16#014A# => return "0000101000001101";
      when 16#014C# => return "0010000000100000";
      when 16#014E# => return "0010000001100111";
      when 16#0150# => return "0010110100100000";
      when 16#0152# => return "0111001000100000";
      when 16#0154# => return "0110111001110101";
      when 16#0156# => return "0110001100100000";
      when 16#0158# => return "0110010001101111";
      when 16#015A# => return "0010000001100101";
      when 16#015C# => return "0111001001100110";
      when 16#015E# => return "0110110101101111";
      when 16#0160# => return "0011000000100000";
      when 16#0162# => return "0011100001111000";
      when 16#0164# => return "0011000000110000";
      when 16#0166# => return "0000110100110000";
      when 16#0168# => return "0000000000001010";
      when 16#016A# => return "0000010100001000";
      when 16#016C# => return "0000000000000010";
      when 16#016E# => return "0000001000001000";
      when 16#0170# => return "0000000110100000";
      when 16#0172# => return "0011110000001000";
      when 16#0174# => return "0110000100000000";
      when 16#0176# => return "0000000100001000";
      when 16#0178# => return "0000000000001010";
      when 16#017A# => return "0000001000001000";
      when 16#017C# => return "1000000000000000";
      when 16#017E# => return "0011000100000000";
      when 16#0180# => return "0011100100000000";
      when 16#0182# => return "0011010000011000";
      when 16#0184# => return "0000100100001000";
      when 16#0186# => return "0000000000000010";
      when 16#0188# => return "0001100110010000";
      when 16#018A# => return "0001000001101010";
      when 16#018C# => return "0100000000000000";
      when 16#018E# => return "0100000100111010";
      when 16#0190# => return "0000000000000001";
      when 16#0192# => return "0000001000001010";
      when 16#0194# => return "0000000110001000";
      when 16#0196# => return "0000000000011000";
      when 16#0198# => return "0011000100000000";
      when 16#019A# => return "0011110000011000";
      when 16#019C# => return "0011010000011000";
      when 16#019E# => return "0000001000011000";
      when 16#01A0# => return "0001010000101000";
      when 16#01A2# => return "0100000000000000";
      when 16#01A4# => return "0000000000011011";
      when 16#01A6# => return "0001010000101000";
      when 16#01A8# => return "0100000000000000";
      when 16#01AA# => return "0000000001011011";
      when 16#01AC# => return "0001010000101000";
      when 16#01AE# => return "0100000000000000";
      when 16#01B0# => return "0000000001001000";
      when 16#01B2# => return "0001010000101000";
      when 16#01B4# => return "0100000000000000";
      when 16#01B6# => return "0000000000011011";
      when 16#01B8# => return "0001010000101000";
      when 16#01BA# => return "0100000000000000";
      when 16#01BC# => return "0000000001011011";
      when 16#01BE# => return "0001010000101000";
      when 16#01C0# => return "0100000000000000";
      when 16#01C2# => return "0000000001001010";
      when 16#01C4# => return "0000001000011000";
      when 16#01C6# => return "0011000100000000";
      when 16#01C8# => return "0011100100000000";
      when 16#01CA# => return "0011010000011000";
      when 16#01CC# => return "0011000100000000";
      when 16#01CE# => return "0011110000011000";
      when 16#01D0# => return "0011010000011000";
      when 16#01D2# => return "0000001000011000";
      when others   => return "0000000000000000";
    end case;
  end function;

end package body;
