LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

package generated is

  function builtin_rom(addr : in std_logic_vector(15 downto 1)) return std_logic_vector;

end package;

package body generated is

  function builtin_rom(addr : in std_logic_vector(15 downto 1)) return std_logic_vector is
  begin
    case to_integer(unsigned(addr & "0")) is
      when 16#0000# => return "0000001000001000";
      when 16#0002# => return "0000000000001010";
      when 16#0004# => return "0000001101010110";
      when 16#0006# => return "0000001100110100";
      when 16#0008# => return "0000001111011110";
      when 16#000A# => return "0011110000001000";
      when 16#000C# => return "0111000000000000";
      when 16#000E# => return "0011010000001000";
      when 16#0010# => return "0111000000000000";
      when 16#0012# => return "0000000100001000";
      when 16#0014# => return "0000000000100100";
      when 16#0016# => return "0000010100001000";
      when 16#0018# => return "0000000000000010";
      when 16#001A# => return "0000001000001000";
      when 16#001C# => return "0000001100110100";
      when 16#001E# => return "0000000000011000";
      when 16#0020# => return "0000001000001000";
      when 16#0022# => return "0000000010001000";
      when 16#0024# => return "0101101100011011";
      when 16#0026# => return "0001101101001000";
      when 16#0028# => return "0100101001011011";
      when 16#002A# => return "0011110100101110";
      when 16#002C# => return "0011110100111101";
      when 16#002E# => return "0011110100111101";
      when 16#0030# => return "0011110100111101";
      when 16#0032# => return "0011110100111101";
      when 16#0034# => return "0011110100111101";
      when 16#0036# => return "0011110100111101";
      when 16#0038# => return "0011110100111101";
      when 16#003A# => return "0011110100111101";
      when 16#003C# => return "0011110100111101";
      when 16#003E# => return "0011110100111101";
      when 16#0040# => return "0011110100111101";
      when 16#0042# => return "0011110100111101";
      when 16#0044# => return "0010111000111101";
      when 16#0046# => return "0000101000001101";
      when 16#0048# => return "0010000001111100";
      when 16#004A# => return "0101001101000001";
      when 16#004C# => return "0100010101001000";
      when 16#004E# => return "0010000001010100";
      when 16#0050# => return "0100111101001000";
      when 16#0052# => return "0100010101001101";
      when 16#0054# => return "0100001100100000";
      when 16#0056# => return "0100110101001111";
      when 16#0058# => return "0101010101010000";
      when 16#005A# => return "0100010101010100";
      when 16#005C# => return "0010000001010010";
      when 16#005E# => return "0100100101000010";
      when 16#0060# => return "0101001101001111";
      when 16#0062# => return "0111110000100000";
      when 16#0064# => return "0000101000001101";
      when 16#0066# => return "0011110100100111";
      when 16#0068# => return "0011110100111101";
      when 16#006A# => return "0011110100111101";
      when 16#006C# => return "0011110100111101";
      when 16#006E# => return "0011110100111101";
      when 16#0070# => return "0011110100111101";
      when 16#0072# => return "0011110100111101";
      when 16#0074# => return "0011110100111101";
      when 16#0076# => return "0011110100111101";
      when 16#0078# => return "0011110100111101";
      when 16#007A# => return "0011110100111101";
      when 16#007C# => return "0011110100111101";
      when 16#007E# => return "0011110100111101";
      when 16#0080# => return "0010011100111101";
      when 16#0082# => return "0000101000001101";
      when 16#0084# => return "0000101000001101";
      when 16#0088# => return "0001010000101000";
      when 16#008A# => return "0100000000000000";
      when 16#008C# => return "0000000000001101";
      when 16#008E# => return "0001010000101000";
      when 16#0090# => return "0100000000000000";
      when 16#0092# => return "0000000000111110";
      when 16#0094# => return "0001010000101000";
      when 16#0096# => return "0100000000000000";
      when 16#0098# => return "0000000000100000";
      when 16#009A# => return "0001010000101000";
      when 16#009C# => return "0100000000000000";
      when 16#009E# => return "0000000000100000";
      when 16#00A0# => return "0001010000101000";
      when 16#00A2# => return "0100000000000000";
      when 16#00A4# => return "0000000000001000";
      when 16#00A6# => return "0001110110001000";
      when 16#00A8# => return "0100000000000000";
      when 16#00AA# => return "0000001001101100";
      when 16#00AC# => return "0000000010100110";
      when 16#00AE# => return "0001010001001000";
      when 16#00B0# => return "0100000000000000";
      when 16#00B2# => return "0100010010110000";
      when 16#00B4# => return "0000000001101000";
      when 16#00B6# => return "0000001001101001";
      when 16#00B8# => return "0000000011011000";
      when 16#00BA# => return "0100010010110000";
      when 16#00BC# => return "0000000001100111";
      when 16#00BE# => return "0000001001101001";
      when 16#00C0# => return "0000000101101110";
      when 16#00C2# => return "0100010010110000";
      when 16#00C4# => return "0000000001111000";
      when 16#00C6# => return "0000001001101001";
      when 16#00C8# => return "0000001101111100";
      when 16#00CA# => return "0100010010110000";
      when 16#00CC# => return "0000000001101100";
      when 16#00CE# => return "0000001001101001";
      when 16#00D0# => return "0000000110000010";
      when 16#00D2# => return "0000000000011000";
      when 16#00D4# => return "0000001000001000";
      when 16#00D6# => return "0000000010001000";
      when 16#00D8# => return "0000000100001000";
      when 16#00DA# => return "0000000011101010";
      when 16#00DC# => return "0000010100001000";
      when 16#00DE# => return "0000000000000010";
      when 16#00E0# => return "0000001000001000";
      when 16#00E2# => return "0000001100110100";
      when 16#00E4# => return "0000000000011000";
      when 16#00E6# => return "0000001000001000";
      when 16#00E8# => return "0000000010001000";
      when 16#00EA# => return "0000101000001101";
      when 16#00EC# => return "0111011001100001";
      when 16#00EE# => return "0110100101100001";
      when 16#00F0# => return "0110000101101100";
      when 16#00F2# => return "0110110001100010";
      when 16#00F4# => return "0010000001100101";
      when 16#00F6# => return "0110111101100011";
      when 16#00F8# => return "0110110101101101";
      when 16#00FA# => return "0110111001100001";
      when 16#00FC# => return "0111001101100100";
      when 16#00FE# => return "0000110100111010";
      when 16#0100# => return "0010000000001010";
      when 16#0102# => return "0110100000100000";
      when 16#0104# => return "0010000000100000";
      when 16#0106# => return "0010000000101101";
      when 16#0108# => return "0110100101100100";
      when 16#010A# => return "0111000001110011";
      when 16#010C# => return "0110000101101100";
      when 16#010E# => return "0010000001111001";
      when 16#0110# => return "0110010101101000";
      when 16#0112# => return "0111000001101100";
      when 16#0114# => return "0000101000001101";
      when 16#0116# => return "0010000000100000";
      when 16#0118# => return "0010000001100111";
      when 16#011A# => return "0010110100100000";
      when 16#011C# => return "0111001000100000";
      when 16#011E# => return "0110111001110101";
      when 16#0120# => return "0110001100100000";
      when 16#0122# => return "0110010001101111";
      when 16#0124# => return "0010000001100101";
      when 16#0126# => return "0111001001100110";
      when 16#0128# => return "0110110101101111";
      when 16#012A# => return "0011000000100000";
      when 16#012C# => return "0011100001111000";
      when 16#012E# => return "0011000000110000";
      when 16#0130# => return "0000110100110000";
      when 16#0132# => return "0010000000001010";
      when 16#0134# => return "0110110000100000";
      when 16#0136# => return "0010000000100000";
      when 16#0138# => return "0010000000101101";
      when 16#013A# => return "0110111101101100";
      when 16#013C# => return "0110010001100001";
      when 16#013E# => return "0010000001110011";
      when 16#0140# => return "0110111001100001";
      when 16#0142# => return "0110100100100000";
      when 16#0144# => return "0110010101101000";
      when 16#0146# => return "0010000001111000";
      when 16#0148# => return "0110100101100110";
      when 16#014A# => return "0110010101101100";
      when 16#014C# => return "0000101000001101";
      when 16#014E# => return "0010000000100000";
      when 16#0150# => return "0010000001111000";
      when 16#0152# => return "0010110100100000";
      when 16#0154# => return "0111010000100000";
      when 16#0156# => return "0111001101100101";
      when 16#0158# => return "0111001101110100";
      when 16#015A# => return "0111001100100000";
      when 16#015C# => return "0111001001100101";
      when 16#015E# => return "0110000101101001";
      when 16#0160# => return "0101111101101100";
      when 16#0162# => return "0110010101110010";
      when 16#0164# => return "0110010001100001";
      when 16#0166# => return "0110110001011111";
      when 16#0168# => return "0110111001101001";
      when 16#016A# => return "0000110101100101";
      when 16#016C# => return "0000000000001010";
      when 16#016E# => return "0000010100001000";
      when 16#0170# => return "0000000000000010";
      when 16#0172# => return "0000001000001000";
      when 16#0174# => return "0000001101010110";
      when 16#0176# => return "0011110000001000";
      when 16#0178# => return "0111000000000000";
      when 16#017A# => return "0000000100001000";
      when 16#017C# => return "0000000000001010";
      when 16#017E# => return "0000001000001000";
      when 16#0180# => return "1000000000000000";
      when 16#0182# => return "0000000100001000";
      when 16#0184# => return "0000001001010010";
      when 16#0186# => return "0000010100001000";
      when 16#0188# => return "0000000000000010";
      when 16#018A# => return "0000001000001000";
      when 16#018C# => return "0000001100110100";
      when 16#018E# => return "0000000000011000";
      when 16#0190# => return "0001110100001000";
      when 16#0192# => return "0100000000000000";
      when 16#0194# => return "0100010010111000";
      when 16#0196# => return "0000000000111010";
      when 16#0198# => return "0000001000001100";
      when 16#019A# => return "0000000110010000";
      when 16#019C# => return "0000000100001000";
      when 16#01A0# => return "0000010100001000";
      when 16#01A2# => return "0000000000000010";
      when 16#01A4# => return "0000001000001000";
      when 16#01A6# => return "0000001001101100";
      when 16#01A8# => return "0000000100001000";
      when 16#01AC# => return "0000010100001000";
      when 16#01AE# => return "0000000000000010";
      when 16#01B0# => return "0000001000001000";
      when 16#01B2# => return "0000001001101100";
      when 16#01B4# => return "0111000100011000";
      when 16#01B6# => return "0000000100001000";
      when 16#01BA# => return "0000010100001000";
      when 16#01BC# => return "0000000000000010";
      when 16#01BE# => return "0000001000001000";
      when 16#01C0# => return "0000001001101100";
      when 16#01C2# => return "0101100101111000";
      when 16#01C4# => return "0000000100001000";
      when 16#01C8# => return "0000010100001000";
      when 16#01CA# => return "0000000000000010";
      when 16#01CC# => return "0000001000001000";
      when 16#01CE# => return "0000001001101100";
      when 16#01D0# => return "0100010010110000";
      when 16#01D4# => return "0000001000001001";
      when 16#01D6# => return "0000000111101010";
      when 16#01D8# => return "0100010010110000";
      when 16#01DA# => return "0000000000000001";
      when 16#01DC# => return "0000001000001001";
      when 16#01DE# => return "0000001000111010";
      when 16#01E0# => return "0000000000011000";
      when 16#01E2# => return "0000000000011000";
      when 16#01E4# => return "0000000000011000";
      when 16#01E6# => return "0000001000001000";
      when 16#01E8# => return "0000000110010000";
      when 16#01EA# => return "0000100110001000";
      when 16#01EC# => return "1111111111111111";
      when 16#01EE# => return "0000001000001001";
      when 16#01F0# => return "0000001000011010";
      when 16#01F2# => return "0000000100001000";
      when 16#01F6# => return "0000010100001000";
      when 16#01F8# => return "0000000000000010";
      when 16#01FA# => return "0000001000001000";
      when 16#01FC# => return "0000001001101100";
      when 16#01FE# => return "0000100100001000";
      when 16#0200# => return "1111111111111110";
      when 16#0202# => return "0100000100110000";
      when 16#0204# => return "0000000000000001";
      when 16#0206# => return "0000110001101000";
      when 16#0208# => return "1111111111111110";
      when 16#020A# => return "0001000001111000";
      when 16#020C# => return "0100010110111000";
      when 16#020E# => return "0000000000000001";
      when 16#0210# => return "0001010000101000";
      when 16#0212# => return "0100000000000000";
      when 16#0214# => return "0000000000101110";
      when 16#0216# => return "0000001000001000";
      when 16#0218# => return "0000000111101110";
      when 16#021A# => return "0000010100001000";
      when 16#021C# => return "0000000000000010";
      when 16#021E# => return "0000001000001000";
      when 16#0220# => return "0000001001101100";
      when 16#0222# => return "0000000000011000";
      when 16#0224# => return "0000000000011000";
      when 16#0226# => return "0000000000011000";
      when 16#0228# => return "0000000000011000";
      when 16#022A# => return "0001010000101000";
      when 16#022C# => return "0100000000000000";
      when 16#022E# => return "0000000000001101";
      when 16#0230# => return "0001010000101000";
      when 16#0232# => return "0100000000000000";
      when 16#0234# => return "0000000000001010";
      when 16#0236# => return "0000001000001000";
      when 16#0238# => return "0000000110010000";
      when 16#023A# => return "0000000100001000";
      when 16#023E# => return "0000010100001000";
      when 16#0240# => return "0000000000000010";
      when 16#0242# => return "0000001000001000";
      when 16#0244# => return "0000001001101100";
      when 16#0246# => return "0000000000011000";
      when 16#0248# => return "0000000000011000";
      when 16#024A# => return "0000000000011000";
      when 16#024C# => return "0000000000011000";
      when 16#024E# => return "0000001000001000";
      when 16#0250# => return "0000000010001000";
      when 16#0252# => return "0000101000001101";
      when 16#0254# => return "0111011101100001";
      when 16#0256# => return "0110100101100001";
      when 16#0258# => return "0110100101110100";
      when 16#025A# => return "0110011101101110";
      when 16#025C# => return "0110100100100000";
      when 16#025E# => return "0110010101101000";
      when 16#0260# => return "0010000001111000";
      when 16#0262# => return "0110100101100110";
      when 16#0264# => return "0110010101101100";
      when 16#0266# => return "0010111000101110";
      when 16#0268# => return "0000110100101110";
      when 16#026A# => return "0000000000001010";
      when 16#026C# => return "0011000100000000";
      when 16#026E# => return "0011100100000000";
      when 16#0270# => return "0011010000011000";
      when 16#0272# => return "0001110100001000";
      when 16#0274# => return "0100000000000000";
      when 16#0276# => return "0110010110011000";
      when 16#0278# => return "0000001001101100";
      when 16#027A# => return "0000001001110010";
      when 16#027C# => return "0100000100111000";
      when 16#027E# => return "0000001010110100";
      when 16#0280# => return "0001100100011000";
      when 16#0282# => return "0110010110011000";
      when 16#0284# => return "0000001001101100";
      when 16#0286# => return "0000001001110010";
      when 16#0288# => return "0111100100011000";
      when 16#028A# => return "0111100100011000";
      when 16#028C# => return "0111100100011000";
      when 16#028E# => return "0111100100011000";
      when 16#0290# => return "0001110100001000";
      when 16#0292# => return "0100000000000000";
      when 16#0294# => return "0110010110011000";
      when 16#0296# => return "0000001001101100";
      when 16#0298# => return "0000001010010000";
      when 16#029A# => return "0100000100111000";
      when 16#029C# => return "0000001010110100";
      when 16#029E# => return "0001100100011000";
      when 16#02A0# => return "0110010110011000";
      when 16#02A2# => return "0000001001101100";
      when 16#02A4# => return "0000001010010000";
      when 16#02A6# => return "0101100101111000";
      when 16#02A8# => return "0000110001101000";
      when 16#02AA# => return "0000000000000010";
      when 16#02AC# => return "0011000100000000";
      when 16#02AE# => return "0011110000011000";
      when 16#02B0# => return "0011010000011000";
      when 16#02B2# => return "0000001000011000";
      when 16#02B4# => return "1111111111111111";
      when 16#02B6# => return "1111111111111111";
      when 16#02B8# => return "1111111111111111";
      when 16#02BA# => return "1111111111111111";
      when 16#02BC# => return "1111111111111111";
      when 16#02BE# => return "1111111111111111";
      when 16#02C0# => return "1111111111111111";
      when 16#02C2# => return "1111111111111111";
      when 16#02C4# => return "1111111111111111";
      when 16#02C6# => return "1111111111111111";
      when 16#02C8# => return "1111111111111111";
      when 16#02CA# => return "1111111111111111";
      when 16#02CC# => return "1111111111111111";
      when 16#02CE# => return "1111111111111111";
      when 16#02D0# => return "1111111111111111";
      when 16#02D2# => return "1111111111111111";
      when 16#02D4# => return "1111111111111111";
      when 16#02D6# => return "1111111111111111";
      when 16#02D8# => return "1111111111111111";
      when 16#02DA# => return "1111111111111111";
      when 16#02DC# => return "1111111111111111";
      when 16#02DE# => return "1111111111111111";
      when 16#02E0# => return "1111111111111111";
      when 16#02E2# => return "1111111111111111";
      when 16#02E4# => return "0000000100000000";
      when 16#02E6# => return "0000001100000010";
      when 16#02E8# => return "0000010100000100";
      when 16#02EA# => return "0000011100000110";
      when 16#02EC# => return "0000100100001000";
      when 16#02EE# => return "1111111111111111";
      when 16#02F0# => return "1111111111111111";
      when 16#02F2# => return "1111111111111111";
      when 16#02F4# => return "0000101011111111";
      when 16#02F6# => return "0000110000001011";
      when 16#02F8# => return "0000111000001101";
      when 16#02FA# => return "1111111100001111";
      when 16#02FC# => return "1111111111111111";
      when 16#02FE# => return "1111111111111111";
      when 16#0300# => return "1111111111111111";
      when 16#0302# => return "1111111111111111";
      when 16#0304# => return "1111111111111111";
      when 16#0306# => return "1111111111111111";
      when 16#0308# => return "1111111111111111";
      when 16#030A# => return "1111111111111111";
      when 16#030C# => return "1111111111111111";
      when 16#030E# => return "1111111111111111";
      when 16#0310# => return "1111111111111111";
      when 16#0312# => return "1111111111111111";
      when 16#0314# => return "0000101011111111";
      when 16#0316# => return "0000110000001011";
      when 16#0318# => return "0000111000001101";
      when 16#031A# => return "1111111100001111";
      when 16#031C# => return "1111111111111111";
      when 16#031E# => return "1111111111111111";
      when 16#0320# => return "1111111111111111";
      when 16#0322# => return "1111111111111111";
      when 16#0324# => return "1111111111111111";
      when 16#0326# => return "1111111111111111";
      when 16#0328# => return "1111111111111111";
      when 16#032A# => return "1111111111111111";
      when 16#032C# => return "1111111111111111";
      when 16#032E# => return "1111111111111111";
      when 16#0330# => return "1111111111111111";
      when 16#0332# => return "1111111111111111";
      when 16#0334# => return "0011000100000000";
      when 16#0336# => return "0011100100000000";
      when 16#0338# => return "0011010000011000";
      when 16#033A# => return "0000100100001000";
      when 16#033C# => return "0000000000000010";
      when 16#033E# => return "0001100110010000";
      when 16#0340# => return "0001000001101010";
      when 16#0342# => return "0100000000000000";
      when 16#0344# => return "0100000100111010";
      when 16#0346# => return "0000000000000001";
      when 16#0348# => return "0000001000001010";
      when 16#034A# => return "0000001100111110";
      when 16#034C# => return "0000000000011000";
      when 16#034E# => return "0011000100000000";
      when 16#0350# => return "0011110000011000";
      when 16#0352# => return "0011010000011000";
      when 16#0354# => return "0000001000011000";
      when 16#0356# => return "0001010000101000";
      when 16#0358# => return "0100000000000000";
      when 16#035A# => return "0000000000011011";
      when 16#035C# => return "0001010000101000";
      when 16#035E# => return "0100000000000000";
      when 16#0360# => return "0000000001011011";
      when 16#0362# => return "0001010000101000";
      when 16#0364# => return "0100000000000000";
      when 16#0366# => return "0000000001001000";
      when 16#0368# => return "0001010000101000";
      when 16#036A# => return "0100000000000000";
      when 16#036C# => return "0000000000011011";
      when 16#036E# => return "0001010000101000";
      when 16#0370# => return "0100000000000000";
      when 16#0372# => return "0000000001011011";
      when 16#0374# => return "0001010000101000";
      when 16#0376# => return "0100000000000000";
      when 16#0378# => return "0000000001001010";
      when 16#037A# => return "0000001000011000";
      when 16#037C# => return "0001010000101000";
      when 16#037E# => return "0100000000000000";
      when 16#0380# => return "0000000000001101";
      when 16#0382# => return "0001010000101000";
      when 16#0384# => return "0100000000000000";
      when 16#0386# => return "0000000000001010";
      when 16#0388# => return "0001010000101000";
      when 16#038A# => return "0100000000000000";
      when 16#038C# => return "0000000000100100";
      when 16#038E# => return "0001010000101000";
      when 16#0390# => return "0100000000000000";
      when 16#0392# => return "0000000000100000";
      when 16#0394# => return "0000000100001000";
      when 16#0396# => return "0000000000100000";
      when 16#0398# => return "0000000100001000";
      when 16#039A# => return "0110000000000000";
      when 16#039C# => return "0000010100001000";
      when 16#039E# => return "0000000000000010";
      when 16#03A0# => return "0000001000001000";
      when 16#03A2# => return "0000001111011110";
      when 16#03A4# => return "0000000000011000";
      when 16#03A6# => return "0000000000011000";
      when 16#03A8# => return "0001010000101000";
      when 16#03AA# => return "0100000000000000";
      when 16#03AC# => return "0000000000001101";
      when 16#03AE# => return "0001010000101000";
      when 16#03B0# => return "0100000000000000";
      when 16#03B2# => return "0000000000001010";
      when 16#03B4# => return "0001010000101000";
      when 16#03B6# => return "0100000000000000";
      when 16#03B8# => return "0000000000111110";
      when 16#03BA# => return "0000000100001000";
      when 16#03BC# => return "0110000000000000";
      when 16#03BE# => return "0000010100001000";
      when 16#03C0# => return "0000000000000010";
      when 16#03C2# => return "0000001000001000";
      when 16#03C4# => return "0000001100110100";
      when 16#03C6# => return "0000000000011000";
      when 16#03C8# => return "0001010000101000";
      when 16#03CA# => return "0100000000000000";
      when 16#03CC# => return "0000000000111100";
      when 16#03CE# => return "0001010000101000";
      when 16#03D0# => return "0100000000000000";
      when 16#03D2# => return "0000000000001101";
      when 16#03D4# => return "0001010000101000";
      when 16#03D6# => return "0100000000000000";
      when 16#03D8# => return "0000000000001010";
      when 16#03DA# => return "0000001000001000";
      when 16#03DC# => return "0000000010001000";
      when 16#03DE# => return "0011000100000000";
      when 16#03E0# => return "0011100100000000";
      when 16#03E2# => return "0011010000011000";
      when 16#03E4# => return "0000000100001000";
      when 16#03E8# => return "0001110110001000";
      when 16#03EA# => return "0100000000000000";
      when 16#03EC# => return "0000001001101100";
      when 16#03EE# => return "0000001111101000";
      when 16#03F0# => return "0100010010110000";
      when 16#03F2# => return "0000000000011011";
      when 16#03F4# => return "0000001000001001";
      when 16#03F6# => return "0000010001110000";
      when 16#03F8# => return "0100010010110000";
      when 16#03FA# => return "0000000000001101";
      when 16#03FC# => return "0000001000001001";
      when 16#03FE# => return "0000010001111000";
      when 16#0400# => return "0100010010110000";
      when 16#0402# => return "0000000001111111";
      when 16#0404# => return "0000001001101001";
      when 16#0406# => return "0000010001000100";
      when 16#0408# => return "0100010010110000";
      when 16#040A# => return "0000000000100000";
      when 16#040C# => return "0000001000001100";
      when 16#040E# => return "0000001111101000";
      when 16#0410# => return "0000100100001000";
      when 16#0412# => return "1111111111111111";
      when 16#0414# => return "0000100100001000";
      when 16#0416# => return "0000000000000011";
      when 16#0418# => return "0100010100111000";
      when 16#041A# => return "0000000000000001";
      when 16#041C# => return "0100010011111000";
      when 16#041E# => return "0000001001101110";
      when 16#0420# => return "0000001111101000";
      when 16#0422# => return "0001000001001000";
      when 16#0424# => return "0100000000000000";
      when 16#0426# => return "0000100100001000";
      when 16#0428# => return "0000000000000010";
      when 16#042A# => return "0000100100001000";
      when 16#042C# => return "1111111111111111";
      when 16#042E# => return "0100000101111000";
      when 16#0430# => return "0001000001111000";
      when 16#0432# => return "0100000100111000";
      when 16#0434# => return "0000000000000001";
      when 16#0436# => return "0000100100001000";
      when 16#0438# => return "0000000000000010";
      when 16#043A# => return "0100000101011000";
      when 16#043C# => return "0001000000111000";
      when 16#0440# => return "0000001000001000";
      when 16#0442# => return "0000001111101000";
      when 16#0444# => return "0100010010110000";
      when 16#0448# => return "0000001000001001";
      when 16#044A# => return "0000001111101000";
      when 16#044C# => return "0100010100111000";
      when 16#044E# => return "0000000000000001";
      when 16#0450# => return "0000100100001000";
      when 16#0452# => return "0000000000000010";
      when 16#0454# => return "0100000101011000";
      when 16#0456# => return "0001000000111000";
      when 16#045A# => return "0001000000101000";
      when 16#045C# => return "0100000000000000";
      when 16#045E# => return "0000000000001000";
      when 16#0460# => return "0001000000101000";
      when 16#0462# => return "0100000000000000";
      when 16#0464# => return "0000000000100000";
      when 16#0466# => return "0001000000101000";
      when 16#0468# => return "0100000000000000";
      when 16#046A# => return "0000000000001000";
      when 16#046C# => return "0000001000001000";
      when 16#046E# => return "0000001111101000";
      when 16#0470# => return "0000100100001000";
      when 16#0472# => return "0000000000000010";
      when 16#0474# => return "0001000000111000";
      when 16#0478# => return "0011000100000000";
      when 16#047A# => return "0011110000011000";
      when 16#047C# => return "0011010000011000";
      when 16#047E# => return "0000001000011000";
      when others   => return "0000000000000000";
    end case;
  end function;

end package body;
