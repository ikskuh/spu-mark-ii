

package SPU_Mark_II_Types is
	TYPE RegisterName IS (
		IR,
		FR,
		IP,
		SP,
		BP
	);		
end package;